module array_gates(output [15:0]o,input [15:0] a, b);
	and(o[0], a[0], b[0]);
	and(o[1], a[1], b[1]);
	and(o[2], a[2], b[2]); 
	and(o[3], a[3], b[3]);
	and(o[4], a[4], b[4]); 
	and(o[5], a[5], b[5]);
	and(o[6], a[6], b[6]); 
	and(o[7], a[7], b[7]); 
	and(o[8], a[8], b[8]); 
	and(o[9], a[9], b[9]); 
	and(o[10], a[10], b[10]); 
	and(o[11], a[11], b[11]); 
	and(o[12], a[12], b[12]); 
	and(o[13], a[13], b[13]); 
	and(o[14], a[14], b[14]); 
	and(o[15], a[15], b[15]); 

endmodule
